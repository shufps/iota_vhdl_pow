entity curlslow is
	port
	(
	);
end curlslow;

architecture behv of curlslow is
begin

end curlslow;
